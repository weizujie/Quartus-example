library verilog;
use verilog.vl_types.all;
entity my_and2 is
    port(
        output_3        : out    vl_logic;
        input1_1        : in     vl_logic;
        input2_2        : in     vl_logic
    );
end my_and2;
