library verilog;
use verilog.vl_types.all;
entity m_faddr_vlg_vec_tst is
end m_faddr_vlg_vec_tst;
