library verilog;
use verilog.vl_types.all;
entity full_addr_vlg_check_tst is
    port(
        CO_7            : in     vl_logic;
        SUM_10          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end full_addr_vlg_check_tst;
