library verilog;
use verilog.vl_types.all;
entity cnt4_to_16_vlg_check_tst is
    port(
        co              : in     vl_logic;
        q               : in     vl_logic_vector(1 downto 0);
        sampler_rx      : in     vl_logic
    );
end cnt4_to_16_vlg_check_tst;
