library verilog;
use verilog.vl_types.all;
entity my_and2_vlg_check_tst is
    port(
        output_3        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end my_and2_vlg_check_tst;
