library verilog;
use verilog.vl_types.all;
entity cnt4_to_16_vlg_vec_tst is
end cnt4_to_16_vlg_vec_tst;
