library verilog;
use verilog.vl_types.all;
entity sled_vlg_vec_tst is
end sled_vlg_vec_tst;
