library verilog;
use verilog.vl_types.all;
entity dled_17990425_vlg_sample_tst is
    port(
        CLK48M          : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end dled_17990425_vlg_sample_tst;
