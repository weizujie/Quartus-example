library verilog;
use verilog.vl_types.all;
entity full_addr_vlg_vec_tst is
end full_addr_vlg_vec_tst;
