library verilog;
use verilog.vl_types.all;
entity half_addr_vlg_vec_tst is
end half_addr_vlg_vec_tst;
