library verilog;
use verilog.vl_types.all;
entity dled_17990425_vlg_vec_tst is
end dled_17990425_vlg_vec_tst;
