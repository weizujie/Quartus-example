library verilog;
use verilog.vl_types.all;
entity my_and2_vlg_vec_tst is
end my_and2_vlg_vec_tst;
